//-------------------------------------------------------------------------------------------------
module sprom
//-------------------------------------------------------------------------------------------------
#
(
	parameter init_file  = "rom8x16K.hex",
	parameter widthad_a = 14,
	parameter width_a = 8
)
(
	input  wire         clock,
	output reg [width_a-1:0] q,
	input  wire[widthad_a-1:0] address
);
//-------------------------------------------------------------------------------------------------

reg[width_a-1:0] d[(2**widthad_a)-1:0];
initial $readmemh(init_file, d, 0);

always @(posedge clock) q<= d[address];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
